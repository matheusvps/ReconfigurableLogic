library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity NiosAndUserHW is
  port(
    clk        : in  std_logic;
    reset_n    : in  std_logic;

    -- Avalon slave (32-bit wide bus typical)
    avs_address    : in  std_logic_vector(1 downto 0); -- vamos mapear 0..3 offsets (00,01,10)
    avs_write      : in  std_logic;
    avs_read       : in  std_logic;
    avs_writedata  : in  std_logic_vector(31 downto 0);
    avs_readdata   : out std_logic_vector(31 downto 0);
    avs_chipselect : in  std_logic
  );
end entity;
architecture rtl of NiosAndUserHW is

  -- registradores internos (8 bits address/data)
  signal reg_addr     : unsigned(9 downto 0) := (others => '0'); -- 10 bits para 1024 endereços
  signal reg_data     : std_logic_vector(7 downto 0) := (others => '0');
  signal reg_control  : std_logic_vector(31 downto 0) := (others => '0');

  -- controle de operações self-clearing
  signal we_mem_pulse : std_logic := '0';
  signal rd_mem_pulse : std_logic := '0';

  -- BRAM signals
  signal bram_addr    : unsigned(9 downto 0);
  signal bram_wren    : std_logic;
  signal bram_din     : std_logic_vector(31 downto 0);
  signal bram_dout    : std_logic_vector(31 downto 0);

  -- readdata combinational
  signal read_data_out : std_logic_vector(31 downto 0);

begin

  -- Decode BRAM signals
  bram_addr <= reg_addr;
  bram_din  <= (31 downto 8 => '0') & reg_data; -- convert 8-bit to 32-bit
  bram_wren <= we_mem_pulse and avs_chipselect;  -- only write if chipselect=1

  -- BRAM instantiation (use the IP generated by Quartus - example port names)
  bram_inst : entity work.bram1024x32
    port map (
      clock    => clk,
      address  => std_logic_vector(bram_addr), -- adjust type to your RAM IP
      wren     => bram_wren,
      data     => bram_din,
      q        => bram_dout
    );

  -- Read path: when rd_mem_pulse and chipselect => drive readdata
  process(clk)
  begin
    if rising_edge(clk) then
      if reset_n = '0' then
        reg_addr <= (others => '0');
        reg_data <= (others => '0');
        reg_control <= (others => '0');
        we_mem_pulse <= '0';
        rd_mem_pulse <= '0';
      else
        -- Avalon write access
        if avs_chipselect = '1' and avs_write = '1' then
          case avs_address is
            when "00" =>
              -- escrever registro de endereço (assumindo escrita em avs_writedata[9:0])
              reg_addr <= unsigned(avs_writedata(9 downto 0));
            when "01" =>
              -- escrever registro de dado (avs_writedata[7:0])
              reg_data <= avs_writedata(7 downto 0);
            when "10" =>
              -- controle: bits por especificação; vamos assumir LSB = WR, next = RD
              reg_control <= avs_writedata;
              if avs_writedata(0) = '1' then  -- WE_MEM bit
                we_mem_pulse <= '1';
              end if;
              if avs_writedata(1) = '1' then  -- RD_MEM bit
                rd_mem_pulse <= '1';
              end if;
            when others =>
              null;
          end case;
        end if;

        -- processar write pulse: realiza gravação e limpa self-clear
        if we_mem_pulse = '1' then
          -- bram_wren é derivado de we_mem_pulse and chipselect -> will write on the same cycle
          we_mem_pulse <= '0'; -- self clear
        end if;

        -- processar read pulse: captura saída BRAM em um registrador de saída
        if rd_mem_pulse = '1' then
          -- le da BRAM (bram_dout já tem o dado lido)
          -- coloca no read_data_out em 32bits (LSB contains 8 bits, resto 0)
          read_data_out <= bram_dout;
          rd_mem_pulse <= '0'; -- self clear
        else
          -- se não houver leitura ativa, mantemos read_data_out inalterado ou z
          null;
        end if;

      end if;
    end if;
  end process;

  -- avs_readdata driven only when avs_chipselect and avs_read
  avs_readdata <= read_data_out when (avs_chipselect = '1' and avs_read = '1') else (others => 'Z'); -- simulation-only tri-state
  -- Nota: alguns ambientes (síntese) não aceitam 'Z' para sinais de saída do módulo; para integração com Avalon
  -- é preferível usar: avs_readdata <= read_data_out when (avs_chipselect='1' and avs_read='1') else (others => '0');

end architecture;
