library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

Entity SlowTotalizer is
	port(
		input : in unsigned(3 downto 0);
		clk   : in std_logic;
		count : out unsigned(2 downto 0)
	);

end entity;

Architecture A_SlowTotalizer of slowTotalizer is
	
	signal i : integer range 0 to 4 := 0;
	signal Internal_Count : unsigned (2 downto 0) := "000";
	signal CurrentInput : unsigned(3 downto 0) := "0000";
	
	begin
		process(clk)
			begin
				if(input = CurrentInput) then
					if (i < 4) then
						if (input(i) = '1') then
							internal_Count <= internal_Count + "001";
						end if;
						i <= i + 1;
					end if;
				else
					currentInput <= input;
					internal_Count <= "000";
					i <= 0;
				end if;
		end process;
		count <= internal_Count;
end architecture;
			
						
					
						
				
				
	

	